module spi_slave(
    input logic spi_clk,    // SPI clk pin
    output logic spi_miso,  // SPI miso pin
    input  logic spi_mosi,  // SPI mosi pin

    input logic clk_sys,    // System clk
    input logic rst,
    output logic [7:0] data_sync,   // Synchronized data
    output logic data_ready_sync    // Valid data in data_sync
);

logic [7:0] shift_reg;
logic [7:0] temp_reg;

logic [7:0] data_pre_sync;
logic data_ready_pre;

logic [2:0] bit_cnt;

logic shift_done;
logic shift_done_dl1;


always_ff @(posedge spi_clk) begin
    if(rst) begin
        shift_reg <= '0;
        bit_cnt <= '0;
        shift_done <= '0;
        shift_done_dl1 <= '0;
    end
    else begin
        shift_reg[7:1] <= shift_reg[6:0];
        shift_reg[0] <= spi_mosi;
        bit_cnt <= bit_cnt + 1;
        if (bit_cnt == 7 ) begin
            temp_reg <= shift_reg;
            shift_done <= 1;
        end
        else begin
            shift_done <= 0;
        end
        shift_done <= shift_done_dl1;
    end
end

// Synchronize data with clk_sys domain
always_ff @(posedge clk_sys) begin
    if (rst) begin
        data_sync <= 0;
        data_pre_sync <= 0;
        data_ready_pre <= 0;
        data_ready_sync <= 0;
    end
    else begin

        // Basic synchronizer on data
        // Generally synchronizing multiple bits of a register requires a more complex synchronization
        // mechanism. This is due to variability in the sampling time in the different registers due
        // to clock skew.
        // In this case it is ok because `temp_reg` is stable for at least an entire clk_sys
        // cycle no matter the alignment of the clocks when data_ready_dl1 is set.
        data_pre_sync <= temp_reg;
        data_sync <= data_pre_sync;

        // Synchronize data ready signal
        data_ready_pre <= shift_done_dl1;
        data_ready_sync <= data_ready_pre;

    end
end

endmodule